magic
tech sky130A
timestamp 1711177935
<< nwell >>
rect -50 -50 250 250
<< nmos >>
rect 95 -200 110 -100
<< pmos >>
rect 95 0 110 200
<< ndiff >>
rect 45 -110 95 -100
rect 45 -190 55 -110
rect 80 -190 95 -110
rect 45 -200 95 -190
rect 110 -110 160 -100
rect 110 -190 125 -110
rect 150 -190 160 -110
rect 110 -200 160 -190
<< pdiff >>
rect 55 190 95 200
rect 55 10 60 190
rect 80 10 95 190
rect 55 0 95 10
rect 110 190 150 200
rect 110 10 125 190
rect 145 10 150 190
rect 110 0 150 10
<< ndiffc >>
rect 55 -190 80 -110
rect 125 -190 150 -110
<< pdiffc >>
rect 60 10 80 190
rect 125 10 145 190
<< poly >>
rect 95 200 110 215
rect 95 -100 110 0
rect 95 -215 110 -200
<< locali >>
rect 55 190 90 200
rect 55 10 60 190
rect 80 10 90 190
rect 55 0 90 10
rect 115 190 150 200
rect 115 10 125 190
rect 145 10 150 190
rect 115 0 150 10
rect 45 -110 90 -100
rect 45 -190 55 -110
rect 80 -190 90 -110
rect 45 -200 90 -190
rect 115 -110 160 -100
rect 115 -190 125 -110
rect 150 -190 160 -110
rect 115 -200 160 -190
<< end >>
